module adderN();
	input [15:0] a;
	input [15:0] b;
	output[16:0] s;

	assign s= a + b;

endmodule